module mux_1_9 #(
    parameter AW = 128
) (
    input   [AW-1 : 0]RDATA         ,
    input   [3    : 0]CTRL_MUX_1_9  ,

    output  [];
);
    
endmodule